/**************************************
* Module: foo
* Date:2014-10-13  
* Author: geisse     
*
* Description: 
***************************************/
module  foo(
    
);
input x;

    bar b(1);
    bar bar(
    	.x(x)
    );

endmodule

