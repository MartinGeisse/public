/**************************************
* Module: bar
* Date:2014-10-13  
* Author: geisse     
*
* Description: 
***************************************/
module  bar(
    input x;
    output z;
);
    z <= x + y;

endmodule

